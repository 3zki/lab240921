* NGSPICE file created from INV3.ext - technology: sky130A

.subckt INV3 A Y VDD GND
X0 a_n60_n1200 A.t0 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.9 pd=6.6 as=0.9 ps=6.6 w=3 l=0.15
X1 a_n60_n1200 A.t1 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=1.98 pd=13.8 as=1.98 ps=13.8 w=6.6 l=0.15
X2 a_605_n1200 a_n60_n1200 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.9 pd=6.6 as=0.9 ps=6.6 w=3 l=0.15
X3 Y.t0 a_605_n1200 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.98 pd=13.8 as=1.98 ps=13.8 w=6.6 l=0.15
X4 a_605_n1200 a_n60_n1200 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.98 pd=13.8 as=1.98 ps=13.8 w=6.6 l=0.15
X5 Y.t1 a_605_n1200 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.9 pd=6.6 as=0.9 ps=6.6 w=3 l=0.15
R0 A.n0 A.t1 1854.09
R1 A.n0 A.t0 546.266
R2 A A.n0 83.556
R3 GND.n7 GND.n6 969.369
R4 GND.n40 GND.n39 908.108
R5 GND.n7 GND.t0 432.432
R6 GND.n40 GND.t2 432.432
R7 GND.n69 GND.t4 432.432
R8 GND.n96 GND.n70 354.577
R9 GND.n2 GND.n1 292.5
R10 GND.n10 GND.n9 292.5
R11 GND.n14 GND.n13 292.5
R12 GND.n19 GND.n18 292.5
R13 GND.n24 GND.n23 292.5
R14 GND.n28 GND.n27 292.5
R15 GND.n32 GND.n31 292.5
R16 GND.n35 GND.n34 292.5
R17 GND.n43 GND.n42 292.5
R18 GND.n47 GND.n46 292.5
R19 GND.n52 GND.n51 292.5
R20 GND.n57 GND.n56 292.5
R21 GND.n61 GND.n60 292.5
R22 GND.n65 GND.n64 292.5
R23 GND.n75 GND.n74 292.5
R24 GND.n93 GND.n91 292.5
R25 GND.n88 GND.n86 292.5
R26 GND.n84 GND.n82 292.5
R27 GND.n79 GND.n77 292.5
R28 GND.n67 GND.n66 292.5
R29 GND.n97 GND.n96 239.365
R30 GND GND.n97 163.617
R31 GND.n8 GND.n7 115.212
R32 GND.n41 GND.n40 115.212
R33 GND.n70 GND.n69 115.212
R34 GND GND.n32 85.487
R35 GND.n54 GND.t3 72
R36 GND.n21 GND.t1 72
R37 GND.n87 GND.t5 72
R38 GND.n9 GND.n8 62.078
R39 GND.n42 GND.n41 62.078
R40 GND.n18 GND.n17 62.077
R41 GND.n51 GND.n50 62.077
R42 GND.n82 GND.n81 62.077
R43 GND.n91 GND.n90 62.077
R44 GND.n74 GND.n73 62.077
R45 GND.n97 GND.n65 54.322
R46 GND.n56 GND.n55 44.535
R47 GND.n34 GND.n33 44.535
R48 GND.n23 GND.n22 44.535
R49 GND.n1 GND.n0 44.535
R50 GND.n61 GND.n59 8.855
R51 GND.n57 GND.n54 8.855
R52 GND.n52 GND.n49 8.855
R53 GND.n47 GND.n45 8.855
R54 GND.n43 GND.n38 8.855
R55 GND.n28 GND.n26 8.855
R56 GND.n24 GND.n21 8.855
R57 GND.n19 GND.n16 8.855
R58 GND.n14 GND.n12 8.855
R59 GND.n10 GND.n5 8.855
R60 GND.n93 GND.n92 8.855
R61 GND.n88 GND.n87 8.855
R62 GND.n84 GND.n83 8.855
R63 GND.n79 GND.n78 8.855
R64 GND.n65 GND.n36 7.595
R65 GND.n32 GND.n3 7.595
R66 GND.n96 GND.n68 7.595
R67 GND.n65 GND.n63 4.845
R68 GND.n32 GND.n30 4.845
R69 GND.n76 GND.n71 4.845
R70 GND.n96 GND.n95 4.845
R71 GND.n62 GND.n61 4.65
R72 GND.n58 GND.n57 4.65
R73 GND.n53 GND.n52 4.65
R74 GND.n48 GND.n47 4.65
R75 GND.n29 GND.n28 4.65
R76 GND.n25 GND.n24 4.65
R77 GND.n20 GND.n19 4.65
R78 GND.n15 GND.n14 4.65
R79 GND.n76 GND.n75 4.65
R80 GND.n94 GND.n93 4.65
R81 GND.n89 GND.n88 4.65
R82 GND.n85 GND.n84 4.65
R83 GND.n80 GND.n79 4.65
R84 GND.n44 GND.n37 2.283
R85 GND.n11 GND.n4 2.283
R86 GND.n44 GND.n43 2.191
R87 GND.n11 GND.n10 2.191
R88 GND.n48 GND.n44 1.451
R89 GND.n15 GND.n11 1.451
R90 GND.n36 GND.n35 0.44
R91 GND.n3 GND.n2 0.44
R92 GND.n75 GND.n72 0.44
R93 GND.n68 GND.n67 0.44
R94 GND.n53 GND.n48 0.195
R95 GND.n58 GND.n53 0.195
R96 GND.n62 GND.n58 0.195
R97 GND.n63 GND.n62 0.195
R98 GND.n20 GND.n15 0.195
R99 GND.n25 GND.n20 0.195
R100 GND.n29 GND.n25 0.195
R101 GND.n30 GND.n29 0.195
R102 GND.n80 GND.n76 0.195
R103 GND.n85 GND.n80 0.195
R104 GND.n89 GND.n85 0.195
R105 GND.n94 GND.n89 0.195
R106 GND.n95 GND.n94 0.195
R107 VDD.n228 VDD.n227 239.59
R108 VDD VDD.n228 153.6
R109 VDD.n227 VDD.n226 127.143
R110 VDD.n151 VDD.n80 127.143
R111 VDD.n75 VDD.n4 127.143
R112 VDD.n194 VDD.t5 118.2
R113 VDD.n120 VDD.t3 118.2
R114 VDD.n44 VDD.t1 118.2
R115 VDD VDD.n75 95.729
R116 VDD.n153 VDD.n152 92.5
R117 VDD.n163 VDD.n161 92.5
R118 VDD.n168 VDD.n166 92.5
R119 VDD.n172 VDD.n170 92.5
R120 VDD.n177 VDD.n175 92.5
R121 VDD.n181 VDD.n179 92.5
R122 VDD.n186 VDD.n184 92.5
R123 VDD.n190 VDD.n188 92.5
R124 VDD.n195 VDD.n193 92.5
R125 VDD.n199 VDD.n197 92.5
R126 VDD.n204 VDD.n202 92.5
R127 VDD.n208 VDD.n206 92.5
R128 VDD.n213 VDD.n211 92.5
R129 VDD.n217 VDD.n215 92.5
R130 VDD.n222 VDD.n220 92.5
R131 VDD.n159 VDD.n157 92.5
R132 VDD.n89 VDD.n87 92.5
R133 VDD.n94 VDD.n92 92.5
R134 VDD.n98 VDD.n96 92.5
R135 VDD.n103 VDD.n101 92.5
R136 VDD.n107 VDD.n105 92.5
R137 VDD.n112 VDD.n110 92.5
R138 VDD.n116 VDD.n114 92.5
R139 VDD.n121 VDD.n119 92.5
R140 VDD.n125 VDD.n123 92.5
R141 VDD.n130 VDD.n128 92.5
R142 VDD.n134 VDD.n132 92.5
R143 VDD.n139 VDD.n137 92.5
R144 VDD.n143 VDD.n141 92.5
R145 VDD.n148 VDD.n146 92.5
R146 VDD.n77 VDD.n76 92.5
R147 VDD.n85 VDD.n83 92.5
R148 VDD.n13 VDD.n11 92.5
R149 VDD.n18 VDD.n16 92.5
R150 VDD.n22 VDD.n20 92.5
R151 VDD.n27 VDD.n25 92.5
R152 VDD.n31 VDD.n29 92.5
R153 VDD.n36 VDD.n34 92.5
R154 VDD.n40 VDD.n38 92.5
R155 VDD.n45 VDD.n43 92.5
R156 VDD.n49 VDD.n47 92.5
R157 VDD.n54 VDD.n52 92.5
R158 VDD.n58 VDD.n56 92.5
R159 VDD.n63 VDD.n61 92.5
R160 VDD.n67 VDD.n65 92.5
R161 VDD.n72 VDD.n70 92.5
R162 VDD.n1 VDD.n0 92.5
R163 VDD.n9 VDD.n7 92.5
R164 VDD.n225 VDD.t4 70.324
R165 VDD.n79 VDD.t2 70.324
R166 VDD.n3 VDD.t0 70.324
R167 VDD.n228 VDD.n151 54.547
R168 VDD.n220 VDD.n219 34.643
R169 VDD.n211 VDD.n210 34.643
R170 VDD.n202 VDD.n201 34.643
R171 VDD.n193 VDD.n192 34.643
R172 VDD.n184 VDD.n183 34.643
R173 VDD.n175 VDD.n174 34.643
R174 VDD.n166 VDD.n165 34.643
R175 VDD.n157 VDD.n156 34.643
R176 VDD.n146 VDD.n145 34.643
R177 VDD.n137 VDD.n136 34.643
R178 VDD.n128 VDD.n127 34.643
R179 VDD.n119 VDD.n118 34.643
R180 VDD.n110 VDD.n109 34.643
R181 VDD.n101 VDD.n100 34.643
R182 VDD.n92 VDD.n91 34.643
R183 VDD.n83 VDD.n82 34.643
R184 VDD.n70 VDD.n69 34.643
R185 VDD.n61 VDD.n60 34.643
R186 VDD.n52 VDD.n51 34.643
R187 VDD.n43 VDD.n42 34.643
R188 VDD.n34 VDD.n33 34.643
R189 VDD.n25 VDD.n24 34.643
R190 VDD.n16 VDD.n15 34.643
R191 VDD.n7 VDD.n6 34.643
R192 VDD.n226 VDD.n225 28.929
R193 VDD.n80 VDD.n79 28.929
R194 VDD.n4 VDD.n3 28.929
R195 VDD.n163 VDD.n162 9.154
R196 VDD.n168 VDD.n167 9.154
R197 VDD.n172 VDD.n171 9.154
R198 VDD.n177 VDD.n176 9.154
R199 VDD.n181 VDD.n180 9.154
R200 VDD.n186 VDD.n185 9.154
R201 VDD.n190 VDD.n189 9.154
R202 VDD.n195 VDD.n194 9.154
R203 VDD.n199 VDD.n198 9.154
R204 VDD.n204 VDD.n203 9.154
R205 VDD.n208 VDD.n207 9.154
R206 VDD.n213 VDD.n212 9.154
R207 VDD.n217 VDD.n216 9.154
R208 VDD.n222 VDD.n221 9.154
R209 VDD.n89 VDD.n88 9.154
R210 VDD.n94 VDD.n93 9.154
R211 VDD.n98 VDD.n97 9.154
R212 VDD.n103 VDD.n102 9.154
R213 VDD.n107 VDD.n106 9.154
R214 VDD.n112 VDD.n111 9.154
R215 VDD.n116 VDD.n115 9.154
R216 VDD.n121 VDD.n120 9.154
R217 VDD.n125 VDD.n124 9.154
R218 VDD.n130 VDD.n129 9.154
R219 VDD.n134 VDD.n133 9.154
R220 VDD.n139 VDD.n138 9.154
R221 VDD.n143 VDD.n142 9.154
R222 VDD.n148 VDD.n147 9.154
R223 VDD.n13 VDD.n12 9.154
R224 VDD.n18 VDD.n17 9.154
R225 VDD.n22 VDD.n21 9.154
R226 VDD.n27 VDD.n26 9.154
R227 VDD.n31 VDD.n30 9.154
R228 VDD.n36 VDD.n35 9.154
R229 VDD.n40 VDD.n39 9.154
R230 VDD.n45 VDD.n44 9.154
R231 VDD.n49 VDD.n48 9.154
R232 VDD.n54 VDD.n53 9.154
R233 VDD.n58 VDD.n57 9.154
R234 VDD.n63 VDD.n62 9.154
R235 VDD.n67 VDD.n66 9.154
R236 VDD.n72 VDD.n71 9.154
R237 VDD.n227 VDD.n154 8.333
R238 VDD.n151 VDD.n78 8.333
R239 VDD.n75 VDD.n2 8.333
R240 VDD.n227 VDD.n224 4.845
R241 VDD.n160 VDD.n155 4.845
R242 VDD.n151 VDD.n150 4.845
R243 VDD.n86 VDD.n81 4.845
R244 VDD.n75 VDD.n74 4.845
R245 VDD.n10 VDD.n5 4.845
R246 VDD.n160 VDD.n159 4.65
R247 VDD.n164 VDD.n163 4.65
R248 VDD.n169 VDD.n168 4.65
R249 VDD.n173 VDD.n172 4.65
R250 VDD.n178 VDD.n177 4.65
R251 VDD.n182 VDD.n181 4.65
R252 VDD.n187 VDD.n186 4.65
R253 VDD.n191 VDD.n190 4.65
R254 VDD.n196 VDD.n195 4.65
R255 VDD.n200 VDD.n199 4.65
R256 VDD.n205 VDD.n204 4.65
R257 VDD.n209 VDD.n208 4.65
R258 VDD.n214 VDD.n213 4.65
R259 VDD.n218 VDD.n217 4.65
R260 VDD.n223 VDD.n222 4.65
R261 VDD.n86 VDD.n85 4.65
R262 VDD.n90 VDD.n89 4.65
R263 VDD.n95 VDD.n94 4.65
R264 VDD.n99 VDD.n98 4.65
R265 VDD.n104 VDD.n103 4.65
R266 VDD.n108 VDD.n107 4.65
R267 VDD.n113 VDD.n112 4.65
R268 VDD.n117 VDD.n116 4.65
R269 VDD.n122 VDD.n121 4.65
R270 VDD.n126 VDD.n125 4.65
R271 VDD.n131 VDD.n130 4.65
R272 VDD.n135 VDD.n134 4.65
R273 VDD.n140 VDD.n139 4.65
R274 VDD.n144 VDD.n143 4.65
R275 VDD.n149 VDD.n148 4.65
R276 VDD.n10 VDD.n9 4.65
R277 VDD.n14 VDD.n13 4.65
R278 VDD.n19 VDD.n18 4.65
R279 VDD.n23 VDD.n22 4.65
R280 VDD.n28 VDD.n27 4.65
R281 VDD.n32 VDD.n31 4.65
R282 VDD.n37 VDD.n36 4.65
R283 VDD.n41 VDD.n40 4.65
R284 VDD.n46 VDD.n45 4.65
R285 VDD.n50 VDD.n49 4.65
R286 VDD.n55 VDD.n54 4.65
R287 VDD.n59 VDD.n58 4.65
R288 VDD.n64 VDD.n63 4.65
R289 VDD.n68 VDD.n67 4.65
R290 VDD.n73 VDD.n72 4.65
R291 VDD.n154 VDD.n153 0.311
R292 VDD.n159 VDD.n158 0.311
R293 VDD.n78 VDD.n77 0.311
R294 VDD.n85 VDD.n84 0.311
R295 VDD.n2 VDD.n1 0.311
R296 VDD.n9 VDD.n8 0.311
R297 VDD.n224 VDD.n223 0.195
R298 VDD.n223 VDD.n218 0.195
R299 VDD.n218 VDD.n214 0.195
R300 VDD.n214 VDD.n209 0.195
R301 VDD.n209 VDD.n205 0.195
R302 VDD.n205 VDD.n200 0.195
R303 VDD.n200 VDD.n196 0.195
R304 VDD.n196 VDD.n191 0.195
R305 VDD.n191 VDD.n187 0.195
R306 VDD.n187 VDD.n182 0.195
R307 VDD.n182 VDD.n178 0.195
R308 VDD.n178 VDD.n173 0.195
R309 VDD.n173 VDD.n169 0.195
R310 VDD.n169 VDD.n164 0.195
R311 VDD.n164 VDD.n160 0.195
R312 VDD.n150 VDD.n149 0.195
R313 VDD.n149 VDD.n144 0.195
R314 VDD.n144 VDD.n140 0.195
R315 VDD.n140 VDD.n135 0.195
R316 VDD.n135 VDD.n131 0.195
R317 VDD.n131 VDD.n126 0.195
R318 VDD.n126 VDD.n122 0.195
R319 VDD.n122 VDD.n117 0.195
R320 VDD.n117 VDD.n113 0.195
R321 VDD.n113 VDD.n108 0.195
R322 VDD.n108 VDD.n104 0.195
R323 VDD.n104 VDD.n99 0.195
R324 VDD.n99 VDD.n95 0.195
R325 VDD.n95 VDD.n90 0.195
R326 VDD.n90 VDD.n86 0.195
R327 VDD.n74 VDD.n73 0.195
R328 VDD.n73 VDD.n68 0.195
R329 VDD.n68 VDD.n64 0.195
R330 VDD.n64 VDD.n59 0.195
R331 VDD.n59 VDD.n55 0.195
R332 VDD.n55 VDD.n50 0.195
R333 VDD.n50 VDD.n46 0.195
R334 VDD.n46 VDD.n41 0.195
R335 VDD.n41 VDD.n37 0.195
R336 VDD.n37 VDD.n32 0.195
R337 VDD.n32 VDD.n28 0.195
R338 VDD.n28 VDD.n23 0.195
R339 VDD.n23 VDD.n19 0.195
R340 VDD.n19 VDD.n14 0.195
R341 VDD.n14 VDD.n10 0.195
R342 Y.n2 Y.t0 129.996
R343 Y.n27 Y.t1 83.228
R344 Y.n19 Y.n18 9.154
R345 Y.n16 Y.n15 9.154
R346 Y.n13 Y.n12 9.154
R347 Y.n10 Y.n9 9.154
R348 Y.n7 Y.n6 9.154
R349 Y.n4 Y.n3 9.154
R350 Y.n1 Y.n0 9.154
R351 Y.n26 Y.n25 8.855
R352 Y.n29 Y.n28 8.855
R353 Y.n23 Y.n22 4.65
R354 Y.n20 Y.n19 4.65
R355 Y.n17 Y.n16 4.65
R356 Y.n14 Y.n13 4.65
R357 Y.n11 Y.n10 4.65
R358 Y.n8 Y.n7 4.65
R359 Y.n5 Y.n4 4.65
R360 Y.n30 Y.n29 4.65
R361 Y.n33 Y.n32 4.65
R362 Y.n27 Y.n26 3.533
R363 Y.n2 Y.n1 3.522
R364 Y.n32 Y.n31 1.272
R365 Y Y.n24 1.005
R366 Y Y.n34 0.885
R367 Y.n22 Y.n21 0.881
R368 Y.n5 Y.n2 0.722
R369 Y.n30 Y.n27 0.711
R370 Y.n8 Y.n5 0.195
R371 Y.n11 Y.n8 0.195
R372 Y.n14 Y.n11 0.195
R373 Y.n17 Y.n14 0.195
R374 Y.n20 Y.n17 0.195
R375 Y.n23 Y.n20 0.195
R376 Y.n24 Y.n23 0.195
R377 Y.n34 Y.n33 0.195
R378 Y.n33 Y.n30 0.195
C0 Y a_605_n1200 0.15fF
C1 Y VDD 1.09fF
C2 VDD A 0.18fF
C3 a_605_n1200 VDD 1.48fF
C4 a_n60_n1200 A 0.14fF
C5 a_n60_n1200 a_605_n1200 0.18fF
C6 a_n60_n1200 VDD 1.50fF
.ends

