* NGSPICE file created from INV12.ext - technology: sky130A

.subckt INV12 A Y VDD GND
X0 GND.t15 a_371_103 a_891_103 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=0.15
X1 GND.t23 a_891_103 Y.t7 GND.t22 sky130_fd_pr__nfet_01v8 ad=0.225 pd=2.1 as=0.1875 ps=1.25 w=0.75 l=0.15
X2 VDD.t7 A.t0 a_371_103 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=2.15 as=0.4125 ps=2.15 w=1.65 l=0.15
X3 Y.t0 a_891_103 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=2.15 as=0.4125 ps=2.15 w=1.65 l=0.15
X4 a_891_103 a_371_103 GND.t13 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=0.15
X5 Y.t6 a_891_103 GND.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=0.15
X6 a_371_103 A.t1 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=2.15 as=0.4125 ps=2.15 w=1.65 l=0.15
X7 VDD.t15 a_371_103 a_891_103 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=2.15 as=0.4125 ps=2.15 w=1.65 l=0.15
X8 VDD.t21 a_891_103 Y.t1 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.9 as=0.4125 ps=2.15 w=1.65 l=0.15
X9 GND.t19 a_891_103 Y.t5 GND.t18 sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=0.15
X10 Y.t3 a_891_103 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=2.15 as=0.4125 ps=2.15 w=1.65 l=0.15
X11 a_891_103 a_371_103 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=2.15 as=0.4125 ps=2.15 w=1.65 l=0.15
X12 VDD.t17 a_891_103 Y.t2 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=2.15 as=0.4125 ps=2.15 w=1.65 l=0.15
X13 GND.t7 A.t2 a_371_103 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=0.15
X14 GND.t11 a_371_103 a_891_103 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=0.15
X15 a_371_103 A.t3 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.225 ps=2.1 w=0.75 l=0.15
X16 a_891_103 a_371_103 GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=0.15
X17 VDD.t3 A.t4 a_371_103 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=2.15 as=0.4125 ps=2.15 w=1.65 l=0.15
X18 VDD.t11 a_371_103 a_891_103 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=2.15 as=0.4125 ps=2.15 w=1.65 l=0.15
X19 GND.t5 A.t5 a_371_103 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=0.15
X20 Y.t4 a_891_103 GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=0.15
X21 a_371_103 A.t6 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=2.15 as=0.495 ps=3.9 w=1.65 l=0.15
X22 a_891_103 a_371_103 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=2.15 as=0.4125 ps=2.15 w=1.65 l=0.15
X23 a_371_103 A.t7 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=0.15
R0 GND GND.t22 999.936
R1 GND.t22 GND.t20 625.136
R2 GND.t20 GND.t18 625.136
R3 GND.t18 GND.t16 625.136
R4 GND.t16 GND.t14 625.136
R5 GND.t14 GND.t12 625.136
R6 GND.t12 GND.t10 625.136
R7 GND.t10 GND.t8 625.136
R8 GND.t8 GND.t4 625.136
R9 GND.t4 GND.t2 625.136
R10 GND.t2 GND.t6 625.136
R11 GND.t6 GND.t0 625.136
R12 GND.n5 GND.t1 297.074
R13 GND.n10 GND.t23 206.723
R14 GND.n9 GND.n0 170.372
R15 GND.n8 GND.n1 170.372
R16 GND.n7 GND.n2 170.372
R17 GND.n6 GND.n3 170.372
R18 GND.n5 GND.n4 170.372
R19 GND.n9 GND.n8 97.882
R20 GND.n8 GND.n7 97.882
R21 GND.n7 GND.n6 97.882
R22 GND.n6 GND.n5 97.882
R23 GND.n10 GND.n9 90.352
R24 GND.n0 GND.t21 40
R25 GND.n0 GND.t19 40
R26 GND.n1 GND.t17 40
R27 GND.n1 GND.t15 40
R28 GND.n2 GND.t13 40
R29 GND.n2 GND.t11 40
R30 GND.n3 GND.t9 40
R31 GND.n3 GND.t5 40
R32 GND.n4 GND.t3 40
R33 GND.n4 GND.t7 40
R34 GND GND.n10 22.588
R35 Y.n4 Y.t7 40
R36 Y.n4 Y.t6 40
R37 Y.n3 Y.t5 40
R38 Y.n3 Y.t4 40
R39 Y.n0 Y.t1 29.848
R40 Y.n0 Y.t3 29.848
R41 Y.n1 Y.t2 29.848
R42 Y.n1 Y.t0 29.848
R43 Y.n5 Y.n3 7.005
R44 Y.n5 Y.n4 6.755
R45 Y.n2 Y.n1 3.572
R46 Y.n2 Y.n0 3.453
R47 Y Y.n2 0.923
R48 Y Y.n5 0.809
R49 A.n0 A.t0 483.762
R50 A.n1 A.t4 434.821
R51 A.n0 A.t1 434.821
R52 A.n2 A.t6 367.585
R53 A.n3 A.t5 339.162
R54 A.n4 A.t2 290.221
R55 A.n3 A.t7 290.221
R56 A.n5 A.t3 222.985
R57 A.n1 A.n0 48.941
R58 A.n2 A.n1 48.941
R59 A.n4 A.n3 48.941
R60 A.n5 A.n4 48.941
R61 A A.n5 5.033
R62 A A.n2 5.033
R63 VDD.n5 VDD.t1 341.185
R64 VDD VDD.t20 340.648
R65 VDD.n10 VDD.t21 250.832
R66 VDD.t20 VDD.t18 224.545
R67 VDD.t18 VDD.t16 224.545
R68 VDD.t16 VDD.t22 224.545
R69 VDD.t22 VDD.t14 224.545
R70 VDD.t14 VDD.t12 224.545
R71 VDD.t12 VDD.t10 224.545
R72 VDD.t10 VDD.t8 224.545
R73 VDD.t8 VDD.t6 224.545
R74 VDD.t6 VDD.t4 224.545
R75 VDD.t4 VDD.t2 224.545
R76 VDD.t2 VDD.t0 224.545
R77 VDD.n5 VDD.n4 167.016
R78 VDD.n6 VDD.n3 167.016
R79 VDD.n7 VDD.n2 167.016
R80 VDD.n8 VDD.n1 167.016
R81 VDD.n9 VDD.n0 167.016
R82 VDD.n9 VDD.n8 97.882
R83 VDD.n8 VDD.n7 97.882
R84 VDD.n7 VDD.n6 97.882
R85 VDD.n6 VDD.n5 97.882
R86 VDD.n10 VDD.n9 90.352
R87 VDD.n4 VDD.t5 29.848
R88 VDD.n4 VDD.t3 29.848
R89 VDD.n3 VDD.t9 29.848
R90 VDD.n3 VDD.t7 29.848
R91 VDD.n2 VDD.t13 29.848
R92 VDD.n2 VDD.t11 29.848
R93 VDD.n1 VDD.t23 29.848
R94 VDD.n1 VDD.t15 29.848
R95 VDD.n0 VDD.t19 29.848
R96 VDD.n0 VDD.t17 29.848
R97 VDD VDD.n10 20.329
C0 VDD Y 0.56fF
C1 a_371_103 a_891_103 0.61fF
C2 VDD a_891_103 1.08fF
C3 VDD a_371_103 1.07fF
C4 Y a_891_103 0.52fF
C5 A a_371_103 0.54fF
C6 VDD A 0.53fF
.ends

