* NGSPICE file created from INV_TEST.ext - technology: sky130A

.subckt INV_TEST A Y VDD GND
X0 VDD.t1 A.t0 Y.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.75 pd=5.6 as=0.75 ps=5.6 w=2.5 l=0.15
X1 GND.t1 A.t1 Y.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
R0 A A.t0 508.934
R1 A A.t1 267.877
R2 Y.n2 Y.t0 129.996
R3 Y Y.t1 43.542
R4 Y.n1 Y.n0 9.154
R5 Y.n5 Y.n4 4.65
R6 Y.n2 Y.n1 3.522
R7 Y Y.n6 0.896
R8 Y.n4 Y.n3 0.881
R9 Y.n5 Y.n2 0.722
R10 Y.n6 Y.n5 0.177
R11 VDD.n2 VDD.t0 150.416
R12 VDD.n9 VDD.t1 118.2
R13 VDD.n20 VDD.n18 92.5
R14 VDD.n10 VDD.n8 92.5
R15 VDD.n16 VDD.n15 92.5
R16 VDD.n5 VDD.n4 92.5
R17 VDD.n4 VDD.n3 34.643
R18 VDD.n8 VDD.n7 34.643
R19 VDD.n15 VDD.n14 34.643
R20 VDD.n3 VDD.n2 28.929
R21 VDD.n5 VDD.n1 9.154
R22 VDD.n10 VDD.n9 9.154
R23 VDD.n20 VDD.n19 9.154
R24 VDD.n17 VDD.n12 4.845
R25 VDD.n11 VDD.n10 4.65
R26 VDD.n21 VDD.n20 4.65
R27 VDD.n17 VDD.n16 4.65
R28 VDD.n6 VDD.n0 2.351
R29 VDD.n6 VDD.n5 2.256
R30 VDD.n11 VDD.n6 1.417
R31 VDD.n16 VDD.n13 0.311
R32 VDD.n21 VDD.n17 0.195
R33 VDD VDD.n21 0.135
R34 VDD VDD.n11 0.059
R35 GND GND.t0 1737.91
R36 GND GND.t1 44.602
C0 VDD Y 0.38fF
C1 A Y 0.15fF
C2 VDD A 0.15fF
.ends

